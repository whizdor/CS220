module encoder_top();
    // Register
    reg [8:0][16:0]a
endmodule